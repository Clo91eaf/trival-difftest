module add (
  input a, 
  input b,
  output c
);
  assign c = 0;
endmodule
